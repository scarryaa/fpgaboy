module memory (
    input logic i_clk,
    input logic i_rst
);

endmodule
