module reg_file (
    input logic i_clk,
    input logic i_rst
);

endmodule
